module ascii_robot

const (
	templates = {
	"0": r"     ___T_     \n    | o o |    \n    |__-__|    \n    /| []|\    \n  ()/|___|\()  \n     |_|_|     \n     /_|_\     ",
	"1": r"    \.===./    \n    | b d |    \n     \_=_/     \n  o==|ooo|==o  \n     |___|     \n    .'._.'.    \n    |_| |_|    ",
	"2": r"     o___o     \n    //0-0\\    \n    |\_-_/|    \n    /|(\)|\    \n   d |___| b   \n    . \_/  .   \n   . .:::.. .  ",
	"3": r"     T___      \n     |[o]|     \n     \_-_/     \n  7--|=0=|--<  \n     |___|     \n     // \\    \n    _\ //_    ",
	"4": r"      )_(      \n     |ooo|     \n     |_#_|     \n .-._/___\_.-. \n ;   \___/   ; \n     (   )     \n    __) (__    ",
	"5": r"     |---|     \n     |6=6|     \n     |_o_|     \n}-. /\--o/\ .-{\n   \" |___| \"   \n      .\".      \n      |_|      ",
	"6": r"     .---.     \n    } - - {    \n     \_0_/     \n   .=[::+]=.   \n ]=' [___] '=[ \n     /| |\     \n    [_] [_]    ",
	"7": r"      Y__      \n    _/o o\_    \n     \_o_/     \n )=o=|L88|=o=( \n )=o=|___|=o=( \n  .  /___\  .  \n. ..:::::::.  .",
	"8": r"     .===.     \n    //d d\\    \n    \_u_//    \n    ,=|x|=.    \n    'c/_\  'c  \n     /| |\     \n    (0) (0)    ",
	"9": r"     _._._     \n    -)o o(-    \n     \_=_/     \n()ooo|\=/|ooo()\n     |___|     \n      |_|      \n     (ooo)     ",
	"a": r"    .=._,=.    \n   ' (q q) `   \n     _)-(_     \n.'c .\"|_|\". n`.\n'--'  /_\  `--'\n    _// \_    \n   /_o| |o_\   ",
	"b": r"      .-.      \n   ._(u u)_.   \n     (_-_)     \n   .=(+++)=.   \no=\"  (___)  \"=o\n     (_|_)     \n     (o|o)     ",
	"c": r"     ,_,_,     \n     \9 9/     \n     /_-_\     \n   ,\"|+  |\".   \n   _\|+__|/_   \n     /  |      \n    _\  |_     ",
	"d": r"     .===./`   \n    /.n n.\    \n    \"\_=_/\"    \n  (m9\:::/\    \n     /___\6    \n     [] []     \n    /:] [:\    ",
	"e": r"      __i      \n     [p q]     \n      ]-[      \n >===]__o[===< \n     [o__]     \n     ]| |[     \n    [_| |_]    ",
	"f": r"   _ _,_,_ _   \n   \( q p )/   \n     \_\"_/     \n  .==|>o<|==:=L\n  '=c|___|     \n     /7 [|     \n   \/7  [|_    ",
}

eyes = {
	"0": "o o",
	"1": "p q",
	"2": "q p",
	"3": "d b",
	"4": "b d",
	"5": "ooo",
	"6": "[o]",
	"7": "9 9",
	"8": "6=6",
	"9": "u u",
	"a": "n n",
	"b": "q q",
	"c": "d d",
	"d": "- -",
	"e": "0 0",
	"f": "O O",
}

mouths = {
	"0": "-",
	"1": "=",
	"2": "o",
	"3": "O",
	"4": "0",
	"5": "#",
	"6": "u",
	"7": "v",
	"8": "n",
	"9": "r",
	"a": "`",
	"b": "^",
	"c": "A",
	"d": "@",
	"e": "e",
	"f": "E",
}

)

